**HP-LQ
*
V1 1 0 AC 1
C11 2 1 1E+04
C12 2 0 1E+04
R2  2 4 1E-10
C3  2 3 1E+03
R4  3 0 2E-10
R5  5 0 2E-10
R6  5 4 2E-10
X1  3 5 4 OPAMP
.AC DEC 200 1.592E+04 1.592E+06
.PLOT AC VDB(6) -60 0
.PLOT AC VP(6) -200 200
.PLOT AC VG(6) 0 3E-06
.TRAN 0.05 10 0
.PLOT TRAN V(6) 0 1.2
.END
*OpAmp Simple Model 1=+in 2=-in 3=Vo
.SUBCKT OPAMP 1 2 3
G0 3 0 1 2 1.E+10
.ENDS OPAMP
*