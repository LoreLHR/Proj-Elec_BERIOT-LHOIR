**LP-HQ
*
V1 1 0 AC 1
R7  1 2 2E-10
C4  3 2 1E+03
R3  3 4 1E+04
C1  4 5 1E+04
R1  4 5 1E+04
R2  5 6 1E+04
R6  6 0 1E+04
X1  2 4 5 OPAMP
X2  6 4 3 OPAMP
.AC DEC 200 1.592E+04 1.592E+06
.PLOT AC VDB(6) -60 0
.PLOT AC VP(6) -200 200
.PLOT AC VG(6) 0 3E-06
.TRAN 0.05 10 0
.PLOT TRAN V(6) 0 1.2
.END
*OpAmp Simple Model 1=+in 2=-in 3=Vo
.SUBCKT OPAMP 1 2 3
G0 3 0 1 2 1.E+10
.ENDS OPAMP
*