**LPN/HPN-MQ                        
*                                   
V1 1 0 AC 1                         
R1  2 1 0.512688                    
R2  2 0 1e+090                      
R5  4 3 2.41167                     
R6  4 0 0.887008                    
R7  1 5 0.234652                    
R8  0 5 0.174266                    
R9  3 5 1                           
C3  2 3 1                           
C4  2 4 1                           
X1  5 4 3 OPAMP                     
.AC DEC 200 1.592E+04 1.592E+06     
.PLOT AC VDB(6) -60 0               
.PLOT AC VP(6) -200 200             
.PLOT AC VG(6) 0 3E-06              
.TRAN 0.05 10 0                     
.PLOT TRAN V(6) 0 1.2               
.END                                
*OpAmp Simple Model 1=+in 2=-in 3=Vo
.SUBCKT OPAMP 1 2 3                 
G0 3 0 1 2 1.E+10                   
.ENDS OPAMP                         
*                                   
