**GP1
*
V1 1 0 AC 1
R1  1 2 1E+03
R2  2 3 1E+04
R3  7 6 1E+04
R4  5 6 1E+03
R5  5 4 1E+04
R7  3 8 1E+04
C6  4 3 1E+04
C8  8 7 1E+04
X1  2 6 5 OPAMP
X2  0 4 3 OPAMP
X3  0 8 7 OPAMP
.AC DEC 200 1.592E+04 1.592E+06
.PLOT AC VDB(6) -60 0
.PLOT AC VP(6) -200 200
.PLOT AC VG(6) 0 3E-06
.TRAN 0.05 10 0
.PLOT TRAN V(6) 0 1.2
.END
*OpAmp Simple Model 1=+in 2=-in 3=Vo
.SUBCKT OPAMP 1 2 3
G0 3 0 1 2 1.E+10
.ENDS OPAMP
*